module mapper_lrn #(
    parameter N_WIDTH = 2,    
    parameter M_WIDTH = 10,   
    parameter E_WIDTH = 6,    
    parameter F_WIDTH = 6,    
    parameter V_WIDTH = 2,    
    parameter ADDR_BUS_WIDTH = 20,    
    parameter DATA_WIDTH     = 16,    
    parameter ROW_MAJOR      = 1     
)(
    input  logic                             core_clk,               
    input  logic                             reset,                  
    input  logic                             start_normalization,    
    input  logic [N_WIDTH-1:0]              dim4,                   
    input  logic [M_WIDTH-1:0]              dim3,                   
    input  logic [E_WIDTH-1:0]              dim2,                   
    input  logic [F_WIDTH-1:0]              dim1,                   
    input  logic [V_WIDTH-1:0]              padding_num,            
    input  logic                             normalized_window,   
    input  logic                             full_flag,              
    input  logic                             div_out_valid,          
    output logic [ADDR_BUS_WIDTH-1:0]        r_addr,                 
    output logic                             r_enable,               
    output logic [ADDR_BUS_WIDTH-1:0]        w_addr,                 
    output logic                             w_enable,               
    output logic                             normalized_layer        
);  

    // Internal signals
    logic [(F_WIDTH + E_WIDTH + M_WIDTH)-1:0] normalized_pixels_count;
    logic [E_WIDTH-1:0] padded_dim2_reg;
    logic [F_WIDTH-1:0] padded_dim1_reg;
    logic [N_WIDTH-1:0] idx4_w, idx4_r;
    logic [M_WIDTH-1:0] idx3_w, idx3_r;
    logic [E_WIDTH-1:0] idx2_w, idx2_r;
    logic [F_WIDTH-1:0] idx1_w, idx1_r;

    // Timing improvement signals
    logic increment_indices_w;
    logic indices_at_max_w;
    logic [3:0] index_stage;
    logic next_idx1_w, next_idx2_w, next_idx3_w, next_idx4_w;
    logic idx1_max, idx2_max, idx3_max, idx4_max;
    logic write_update_valid;

    // Address computation signals
    logic [F_WIDTH + E_WIDTH-1:0] r_temp_1, r_temp_2; 
    logic [F_WIDTH + E_WIDTH + M_WIDTH-1:0] r_temp_3, r_temp_4; 
    logic [F_WIDTH + E_WIDTH + M_WIDTH + N_WIDTH-1:0] r_temp_5;

    logic [V_WIDTH + E_WIDTH-1:0] w_temp_1; 
    logic [V_WIDTH + F_WIDTH-1:0] w_temp_2; 
    logic [E_WIDTH + V_WIDTH + F_WIDTH-1:0] w_temp_3; 
    logic [F_WIDTH + E_WIDTH-1:0] w_temp_4; 
    logic [F_WIDTH + E_WIDTH + M_WIDTH-1:0] w_temp_5, w_temp_6; 
    logic [F_WIDTH + E_WIDTH + M_WIDTH + N_WIDTH-1:0] w_temp_7;

    // Pipeline registers for address calculation
    logic [ADDR_BUS_WIDTH-1:0] w_sum1, w_sum2, w_sum3;
    logic [ADDR_BUS_WIDTH-1:0] w_addr_temp, r_addr_temp;
    logic [ADDR_BUS_WIDTH-1:0] aligned_w_addr;

    // Padding calculation with registered outputs
    always_ff @(posedge core_clk or posedge reset) begin
        if (reset) begin
            padded_dim2_reg <= '0;
            padded_dim1_reg <= '0;
        end else begin
            padded_dim2_reg <= dim2 + (padding_num << 1);
            padded_dim1_reg <= dim1 + (padding_num << 1);
        end
    end

    // Register comparison results
    always_ff @(posedge core_clk or posedge reset) begin
        if (reset) begin
            idx1_max <= 1'b0;
            idx2_max <= 1'b0;
            idx3_max <= 1'b0;
            idx4_max <= 1'b0;
        end else begin
            idx1_max <= (idx1_w == dim1-1);
            idx2_max <= (idx2_w == dim2-1);
            idx3_max <= (idx3_w == dim3-1);
            idx4_max <= (idx4_w == dim4-1);
        end
    end

    // Write update synchronization
    always_ff @(posedge core_clk or posedge reset) begin
        if (reset) begin
            write_update_valid <= 1'b0;
        end else begin
            write_update_valid <= w_enable && !normalized_layer;
        end
    end

// Separate block for index calculations
    always_ff @(posedge core_clk or posedge reset) begin
        if (reset) begin
            next_idx1_w <= 1'b0;
            next_idx2_w <= 1'b0;
            next_idx3_w <= 1'b0;
            next_idx4_w <= 1'b0;
            index_stage <= 4'b0;
        end else if (increment_indices_w) begin
            case (index_stage)
                4'd0: begin
                    next_idx4_w <= idx4_max ? '0 : idx4_w + 1'b1;
                    index_stage <= 4'd1;
                end
                4'd1: begin
                    if (idx4_max) begin
                        next_idx3_w <= idx3_max ? '0 : idx3_w + 1'b1;
                    end
                    index_stage <= 4'd2;
                end
                4'd2: begin
                    if (idx4_max && idx3_max) begin
                        next_idx2_w <= idx2_max ? '0 : idx2_w + 1'b1;
                    end
                    index_stage <= 4'd3;
                end
                4'd3: begin
                    if (idx4_max && idx3_max && idx2_max) begin
                        next_idx1_w <= idx1_max ? '0 : idx1_w + 1'b1;
                    end
                    index_stage <= 4'd0;
                end
                default: index_stage <= 4'd0;
            endcase
        end
    end

    // Address computation instantiations
    unsigned_wallace_tree_multiplier #(.in1_width(F_WIDTH),.in2_width(E_WIDTH)) R_1(
        .in1(idx1_r),
        .in2(dim2),
        .out(r_temp_1)
    );

    unsigned_wallace_tree_multiplier #(.in1_width(F_WIDTH),.in2_width(E_WIDTH)) R_2(
        .in1(dim1),
        .in2(dim2),
        .out(r_temp_2)
    );

    unsigned_wallace_tree_multiplier #(.in1_width(F_WIDTH + E_WIDTH),.in2_width(M_WIDTH)) R_3(
        .in1(r_temp_2),
        .in2(idx3_r),
        .out(r_temp_3)
    );

    unsigned_wallace_tree_multiplier #(.in1_width(F_WIDTH + E_WIDTH),.in2_width(M_WIDTH)) R_4(
        .in1(r_temp_2),
        .in2(dim3),
        .out(r_temp_4)
    );

    unsigned_wallace_tree_multiplier #(.in1_width(F_WIDTH + E_WIDTH + M_WIDTH),.in2_width(N_WIDTH)) R_5(
        .in1(r_temp_4),
        .in2(idx4_r),
        .out(r_temp_5)
    );

    // Modified CLA instantiations
    cla #(.width(V_WIDTH + E_WIDTH)) W_1(
        .x({{(E_WIDTH){1'b0}}, padding_num}),
        .y({{(V_WIDTH){1'b0}}, idx2_w}),
        .sum(w_temp_1)
    );

    cla #(.width(V_WIDTH + F_WIDTH)) W_2(
        .x({{(F_WIDTH){1'b0}}, padding_num}),
        .y({{(V_WIDTH){1'b0}}, idx1_w}),
        .sum(w_temp_2)
    );

    unsigned_wallace_tree_multiplier #(.in1_width(E_WIDTH),.in2_width(V_WIDTH + F_WIDTH)) W_3(
        .in1(padded_dim2_reg),
        .in2(w_temp_2),
        .out(w_temp_3)
    );

    unsigned_wallace_tree_multiplier #(.in1_width(F_WIDTH),.in2_width(E_WIDTH)) W_4(
        .in1(padded_dim1_reg),
        .in2(padded_dim2_reg),
        .out(w_temp_4)
    );

    unsigned_wallace_tree_multiplier #(.in1_width(F_WIDTH + E_WIDTH),.in2_width(M_WIDTH)) W_5(
        .in1(w_temp_4),
        .in2(idx3_w),
        .out(w_temp_5)
    );
 
    unsigned_wallace_tree_multiplier #(.in1_width(F_WIDTH + E_WIDTH),.in2_width(M_WIDTH)) W_6(
        .in1(w_temp_4),
        .in2(dim3),
        .out(w_temp_6)
    );
   
    unsigned_wallace_tree_multiplier #(.in1_width(F_WIDTH + E_WIDTH + M_WIDTH),.in2_width(N_WIDTH)) W_7(
        .in1(w_temp_6),
        .in2(idx4_w),
        .out(w_temp_7)
    );

    // Pipeline stages for address calculation
    always_ff @(posedge core_clk or posedge reset) begin
        if (reset) begin
            w_sum1 <= '0;
            w_sum2 <= '0;
            w_sum3 <= '0;
            w_addr_temp <= '0;
            r_addr_temp <= '0;
            aligned_w_addr <= '0;
        end else begin
            // Pipeline stages for write address
            w_sum1 <= w_temp_7 + w_temp_5;
            w_sum2 <= w_temp_3 + w_temp_1;
            w_sum3 <= w_sum1 + w_sum2;
            w_addr_temp <= w_sum3;
            aligned_w_addr <= {w_addr_temp[ADDR_BUS_WIDTH-1:2], 2'b00};
            
            // Read address calculation
            r_addr_temp <= r_temp_5 + r_temp_3 + r_temp_1 + idx2_r;
        end
    end

    // Address assignments
    assign w_addr = aligned_w_addr;
    assign r_addr = r_addr_temp;

    // State definitions
    typedef enum logic [2:0] {
        IDLE      = 3'b000,
        WAIT      = 3'b001,
        READ      = 3'b010,
        PROCESS   = 3'b011,
        WRITE     = 3'b100
    } state_t;
    
    (* fsm_encoding = "gray" *)
    state_t current_state, next_state;

    // State Memory
    always_ff @(posedge core_clk or posedge reset) begin
        if (reset)
            current_state <= IDLE;
        else 
            current_state <= next_state;
    end  

    // Next State Logic
    always_comb begin
        next_state = current_state; // Default assignment
        case(current_state) 
            IDLE: begin
                next_state = start_normalization ? READ : IDLE;
            end
            
            READ: begin 
                if(full_flag) begin
                    next_state = PROCESS; 
                end else begin
                    next_state = READ; 
                end
            end 

            PROCESS: begin
                if(normalized_layer) begin
                    next_state = IDLE; 
                end
                else if(div_out_valid) begin
                    next_state = WRITE;         
                end else if (normalized_window) begin
                    next_state = WAIT;
                end else begin
                    next_state = PROCESS;       
                end
            end

            WRITE: begin
                if(!normalized_window) begin
                    next_state = PROCESS;           
                end
                else begin
                    next_state = WRITE;             
                end
            end 

            WAIT: begin
                next_state = READ; 
            end

            default: next_state = IDLE;
        endcase 
    end

    // Output Logic with explicit defaults
    always_ff @(posedge core_clk or posedge reset) begin
        if (reset) begin
            idx4_r <= '0;
            idx3_r <= '0;
            idx2_r <= '0;
            idx1_r <= '0;
            idx4_w <= '0;
            idx3_w <= '0;
            idx2_w <= '0;
            idx1_w <= '0;
            w_enable <= 1'b0;
            r_enable <= 1'b0;
            normalized_pixels_count <= '0;
            normalized_layer <= 1'b0;
            increment_indices_w <= 1'b0;
        end
        else begin           
            // Default assignments to prevent latches
            w_enable <= 1'b0;
            r_enable <= 1'b0;
            increment_indices_w <= 1'b0;
            
            case (current_state)
                IDLE: begin
                    idx4_r <= '0;
                    idx3_r <= '0;
                    idx2_r <= '0;
                    idx1_r <= '0;
                    idx4_w <= '0;
                    idx3_w <= '0;
                    idx2_w <= '0;
                    idx1_w <= '0;
                    normalized_pixels_count <= '0;
                    normalized_layer <= 1'b0;

                    if(next_state == READ) r_enable <= 1'b1;
                end

                READ: begin
                    w_enable <= 1'b0;
                    if (idx3_r == dim3-1) r_enable <= 1'b0;
                    else r_enable <= 1'b1;
                    
                    if(r_enable) begin
                        if (idx4_r == dim4-1) begin
                            idx4_r <= '0;
                            if (idx3_r == dim3-1) begin
                                idx3_r <= '0;
                                if (idx2_r == dim2-1) begin
                                    idx2_r <= '0;
                                    if (idx1_r == dim1-1) begin
                                        idx1_r <= '0;
                                    end
                                    else begin
                                        idx1_r <= idx1_r + 1'b1;
                                    end
                                end
                                else idx2_r <= idx2_r + 1'b1;
                            end
                            else idx3_r <= idx3_r + 1'b1;
                        end
                        else idx4_r <= idx4_r + 1'b1;
                    end
                end

                PROCESS: begin
                    r_enable <= 1'b0;
                    normalized_layer <= 1'b0; 
                    if(div_out_valid) begin
                        w_enable <= 1'b1;
                        normalized_pixels_count <= normalized_pixels_count + 1'b1;
                    end
                end

                WRITE: begin
                    w_enable <= 1'b0;
                    r_enable <= 1'b0;
                    
                    if (normalized_pixels_count == dim1 * dim2 * dim3 * dim4) begin
                        normalized_pixels_count <= '0;
                        normalized_layer <= 1'b1;
                    end

                    if (write_update_valid) begin
                        increment_indices_w <= 1'b1;
                        idx4_w <= next_idx4_w;
                        idx3_w <= next_idx3_w;
                        idx2_w <= next_idx2_w;
                        idx1_w <= next_idx1_w;
                    end else begin
                        increment_indices_w <= 1'b0;
                    end
                end

                WAIT: begin
                    if(next_state == IDLE) r_enable <= 1'b0;
                    else                   r_enable <= 1'b1;
                    normalized_layer <= 1'b0;
                    increment_indices_w <= 1'b0;
                end

                default: begin
                    w_enable <= 1'b0;
                    r_enable <= 1'b0;
                    increment_indices_w <= 1'b0;
                end
            endcase 
        end
    end

endmodule
